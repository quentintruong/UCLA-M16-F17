// EEM16 - Logic Design
// Design Assignment #2 - Problem #2.2
// constants2_2.vh
// Verilog template

`ifndef _constants2_2_vh_
`define _constants2_2_vh_

`define THRESHOLD 2

// These three commands must exist
// Add additional commands if necessary
// Be sure to update the width if required
`define CMD_WIDTH 2
`define CMD_CLEAR (`CMD_WIDTH'd0)
`define CMD_LOAD (`CMD_WIDTH'd1)
`define CMD_HOLD (`CMD_WIDTH'd2)

`endif
